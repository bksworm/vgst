module gst


struct Bus  {
mut:
	b &C.GstBus
}