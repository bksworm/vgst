module gst 

fn test_gst(){
	
}
